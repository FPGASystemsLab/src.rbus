//=============================================================================================
//    Main contributors                         
//      - Jakub Siast         <mailto:jakubsiast@gmail.com>
//=============================================================================================
`default_nettype none
//---------------------------------------------------------------------------------------------
`timescale 1ns / 1ns                            
//=============================================================================================
module eco32_ethernet_ptr   
#
(
 parameter  BUFF_ADDR_WIDTH = 'd8
)   
(                                                                                                                               
input  wire                           clk, 
input  wire                           rst,      
                                   
input  wire                           pa_i_stb,  
input  wire                           pa_i_wen,  
input  wire                    [35:0] pa_i_data,  
input  wire     [BUFF_ADDR_WIDTH-2:0] pa_i_addr, 

output wire                           pa_o_stb,  
output wire                    [35:0] pa_o_data,  

input  wire                           pb_i_stb,  
input  wire                           pb_i_wen,  
input  wire                    [35:0] pb_i_data,  
input  wire     [BUFF_ADDR_WIDTH-2:0] pb_i_addr,  

output wire                           pb_o_stb,  
output wire                    [35:0] pb_o_data
);                                         
//=============================================================================================
// parameters
//============================================================================================= 
localparam          _AW                 =                                    (BUFF_ADDR_WIDTH);
localparam          _MS                 =                                 1<<(BUFF_ADDR_WIDTH);       
//=============================================================================================
// variables                               
//============================================================================================= 
(*ramstyle="no_rw_check"*)  reg     [   35:0]   mem [_MS-1:0];
                            reg     [_AW-1:0]   mem_ptr_a;  
                            reg     [_AW-1:0]   mem_ptr_b;  
//----------------------------------------------------------------------------------------------
                            reg                 pa0_stb;                    
                            reg                 pa1_stb;                    
                            reg        [35:0]   pa1_data;                   
//----------------------------------------------------------------------------------------------
                            reg                 pb0_stb;                    
                            reg                 pb1_stb;                    
                            reg        [35:0]   pb1_data;                   
//==============================================================================================
// port A
//==============================================================================================
wire    [_AW-1:0] pa_x_addr         =                                          {1'b0,pa_i_addr};
//----------------------------------------------------------------------------------------------
always@(posedge clk)
     begin
        if(pa_i_wen) mem[pa_x_addr] <= pa_i_data;
        mem_ptr_a                   <= pa_x_addr;
     end
//---------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)  
    begin    
        pa0_stb                     <=                                                      'd0;
    end
 else 
    begin    
        pa0_stb                     <=                                    !pa_i_wen && pa_i_stb;
    end
//----------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)  
    begin                                                                            
        pa1_stb                     <=                                                      'd0;
        pa1_data                    <=                                                      'd0;
    end
 else 
    begin    
        pa1_stb                     <=                                                  pa0_stb;
        pa1_data                    <=                                           mem[mem_ptr_a];
    end
//----------------------------------------------------------------------------------------------
assign  pa_o_stb                    =                                                   pa1_stb;
assign  pa_o_data                   =                                                  pa1_data;
//==============================================================================================
// port B
//==============================================================================================
wire    [_AW-1:0] pb_x_addr         =                                          {1'b1,pb_i_addr};
//----------------------------------------------------------------------------------------------
always@(posedge clk)
     begin                                                                                                                                                            
        if(pb_i_wen) mem[pb_x_addr] <= pb_i_data;
        mem_ptr_b                   <= pb_x_addr;
     end
//----------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)  
    begin    
        pb0_stb                     <=                                                      'd0;
    end
 else 
    begin    
        pb0_stb                     <=                                    !pb_i_wen && pb_i_stb;
    end
//----------------------------------------------------------------------------------------------
always@(posedge clk or posedge rst)
 if(rst)  
    begin                                                                            
        pb1_stb                     <=                                                      'd0;
        pb1_data                    <=                                                      'd0;
    end
 else 
    begin    
        pb1_stb                     <=                                                  pb0_stb;
        pb1_data                    <=                                           mem[mem_ptr_b];
    end
//----------------------------------------------------------------------------------------------
assign  pb_o_stb                    =                                                   pb1_stb;
assign  pb_o_data                   =                                                  pb1_data;
//============================================================================================= 
endmodule
